`timescale 1ns / 1ps`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/23/2024 12:24:46 AM
// Design Name: 
// Module Name: controller_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

static int arar[16900]= '{183,183,183,182,180,179,184,185,181,185,188,185,180,178,176,175,179,185,187,191,193,194,196,198,200,201,204,207,209,210,210,211,212,209,211,211,210,210,213,215,216,215,216,218,219,220,220,219,218,219,217,215,215,216,217,216,215,214,215,214,212,211,211,212,211,212,212,211,210,211,212,211,210,211,210,209,209,209,208,208,208,210,208,206,206,206,206,205,205,206,204,203,203,202,200,199,199,200,197,198,197,196,195,192,193,195,193,192,193,193,192,190,189,190,188,190,191,190,188,185,186,185,186,187,189,190,190,190,189,189,183,183,183,182,180,179,184,185,181,185,188,185,180,178,176,175,179,185,187,191,193,194,196,198,200,201,204,207,209,210,210,211,212,209,211,211,210,210,213,215,216,215,216,218,219,220,220,219,218,219,217,215,215,216,217,216,215,214,215,214,212,211,211,212,211,212,212,211,210,211,212,211,210,211,210,209,209,209,208,208,208,210,208,206,206,206,206,205,205,206,204,203,203,202,200,199,199,200,197,198,197,196,195,192,193,195,193,192,193,193,192,190,189,190,188,190,191,190,188,185,186,185,186,187,189,190,190,190,189,189,186,186,185,183,181,180,184,187,185,186,184,177,173,173,176,184,195,192,193,196,197,198,200,203,205,208,210,212,214,214,214,214,215,215,217,217,216,216,217,218,219,219,219,220,220,221,221,220,219,218,217,215,215,215,216,215,214,214,214,214,212,212,212,212,211,212,213,213,212,211,211,211,211,210,209,209,209,209,208,208,209,211,209,207,206,206,206,206,207,205,204,203,203,202,201,200,200,199,196,197,194,193,193,192,195,192,191,191,192,192,190,190,191,190,188,190,190,191,190,187,187,188,190,192,193,194,194,195,196,196,185,185,183,182,180,178,180,183,183,184,173,166,174,188,193,192,193,195,197,200,202,203,205,208,210,211,212,213,214,214,214,214,214,216,217,217,216,216,217,217,217,215,215,215,215,215,216,216,215,217,216,215,215,215,215,214,214,215,215,214,213,213,214,213,211,212,213,214,213,211,211,211,211,209,208,208,208,208,208,208,208,209,207,206,206,207,206,206,206,205,204,203,202,202,201,200,200,199,197,197,194,193,194,193,196,191,192,193,194,192,190,191,193,193,191,191,190,191,191,187,186,186,189,192,194,195,195,196,196,196,188,188,185,184,184,182,181,181,181,170,174,182,192,194,192,193,200,198,201,204,206,208,208,209,209,208,209,209,210,210,210,210,210,211,211,211,212,212,213,212,212,212,213,213,213,213,214,215,214,215,215,215,215,214,214,214,214,214,215,215,214,214,215,214,212,213,213,213,212,211,211,211,211,210,209,209,209,209,208,208,208,207,206,207,208,208,207,206,205,206,205,204,203,202,201,200,199,199,197,198,197,197,197,194,195,193,194,195,195,193,191,191,193,195,192,192,190,191,193,188,186,186,188,192,195,197,196,196,195,195,191,191,186,185,187,187,184,183,183,183,183,187,193,195,197,199,201,204,206,208,209,208,208,207,207,207,207,207,208,209,209,209,209,209,208,209,210,211,211,211,210,211,212,213,213,214,215,215,215,214,214,214,214,213,213,214,214,213,215,215,214,214,214,214,213,214,213,212,211,211,211,211,210,210,210,209,209,209,208,207,207,207,206,207,207,207,206,206,206,205,205,204,202,202,201,201,200,199,197,198,197,198,198,194,193,194,193,194,194,193,192,192,193,193,191,191,190,192,195,191,189,188,188,190,192,194,195,195,194,194,190,190,185,184,187,188,188,188,187,192,193,195,195,195,198,201,201,203,204,205,205,205,206,206,207,209,209,209,209,210,210,210,209,209,209,209,211,212,211,211,211,211,212,213,213,214,214,214,214,215,215,215,214,214,214,214,214,214,216,216,215,214,214,214,214,213,213,211,210,211,211,211,210,207,207,206,207,206,205,204,205,207,205,204,204,204,204,204,205,203,203,202,201,201,201,201,200,199,196,197,195,196,198,194,193,194,193,192,194,194,194,193,193,193,191,191,190,192,194,191,191,190,188,187,187,190,192,193,193,193,192,192,188,188,191,192,193,194,194,195,195,198,200,198,199,200,198,199,200,201,202,203,204,205,206,208,209,209,210,210,210,209,209,209,209,209,211,211,211,211,212,212,214,215,215,215,215,215,215,215,215,215,215,215,215,214,213,214,215,215,214,213,214,214,213,213,213,213,212,212,212,211,210,207,207,206,207,206,205,205,205,207,205,204,204,203,203,204,205,203,203,202,201,201,202,202,200,198,197,198,196,196,198,196,195,196,194,193,194,195,195,194,194,194,191,191,191,191,192,190,191,192,191,189,189,190,192,194,195,195,192,192,190,191,194,194,194,194,194,198,195,197,198,197,199,201,199,199,200,202,203,204,204,204,204,207,207,208,209,209,209,209,209,209,208,209,211,211,211,212,213,212,213,214,214,214,214,215,215,215,215,215,215,215,214,212,211,213,213,212,211,212,213,213,211,212,213,214,214,213,212,211,211,211,210,210,211,211,210,210,210,208,208,208,208,208,206,206,206,205,206,205,203,203,204,204,202,198,198,201,199,199,201,198,198,198,195,194,195,195,194,193,193,193,189,190,191,191,191,190,194,190,190,190,191,191,192,193,193,193,193,193,193,192,191,192,192,193,196,194,196,197,195,196,199,201,200,201,201,203,204,205,205,204,203,206,207,208,209,209,209,209,208,209,210,210,210,210,211,212,214,212,214,215,216,216,216,216,216,216,216,217,216,214,212,212,213,214,214,213,213,214,214,213,213,213,214,214,212,211,212,212,212,212,211,211,210,210,209,210,211,209,208,208,210,210,208,207,208,207,206,205,205,205,205,205,205,203,201,200,200,200,200,198,196,196,195,198,195,197,194,195,194,196,191,191,190,187,189,193,190,191,192,191,194,193,199,197,192,192,192,192,193,192,191,192,192,192,195,194,195,196,196,197,199,200,200,202,203,204,205,205,205,205,205,205,206,207,208,209,209,209,209,211,211,212,211,211,212,214,215,215,216,217,217,217,217,217,217,217,218,219,218,216,215,215,216,216,215,215,215,216,216,215,215,213,214,214,212,211,212,212,212,212,211,211,211,211,211,211,212,210,209,209,209,210,209,208,208,207,206,205,204,204,205,205,205,204,202,201,202,200,197,196,198,199,198,199,196,198,195,197,196,197,194,193,193,191,191,193,190,181,187,194,194,192,194,198,198,198,191,191,192,191,191,192,192,192,194,195,195,197,198,199,200,201,202,203,203,204,204,205,206,207,207,206,207,208,209,210,211,211,211,213,213,213,213,213,214,215,217,217,217,218,217,217,217,218,217,218,219,219,219,218,217,217,218,217,217,217,217,217,217,217,217,214,214,214,214,213,213,214,213,212,211,211,211,212,211,212,212,211,210,209,209,209,209,208,209,208,207,206,205,205,205,205,205,204,202,203,204,201,197,197,201,202,200,201,198,199,197,199,199,198,198,197,197,197,196,195,194,191,193,199,197,197,194,197,194,194,190,190,192,191,191,192,192,192,194,197,196,198,200,201,200,202,204,204,204,205,205,206,207,208,209,209,209,210,211,212,212,212,213,214,214,215,214,215,215,216,218,218,218,218,217,217,218,219,219,219,219,220,220,219,218,218,219,218,218,218,218,217,217,217,217,215,215,215,215,215,215,215,215,214,213,212,212,211,211,210,211,210,210,209,209,209,209,208,208,208,208,207,206,206,206,205,204,204,203,204,204,202,199,200,203,202,201,201,199,199,199,200,200,198,200,199,199,201,200,198,198,200,198,200,200,202,201,200,195,195,191,191,193,193,191,193,193,194,195,199,198,199,201,202,201,202,205,205,205,207,207,208,208,209,210,210,211,212,212,213,214,214,214,215,215,215,215,215,216,217,218,218,219,218,218,219,220,220,220,220,220,221,221,220,220,219,219,219,219,219,218,218,217,217,217,216,216,216,216,216,216,216,216,216,214,213,213,212,211,210,210,211,211,210,210,210,210,209,208,208,208,207,207,207,206,204,203,203,204,205,203,202,202,203,203,202,202,200,201,200,200,199,200,199,199,199,199,201,200,199,200,200,199,200,203,200,201,200,199,199,193,193,195,195,193,194,195,196,197,200,199,199,201,202,201,202,205,205,206,207,208,209,209,210,210,210,211,212,213,214,214,215,215,215,215,215,215,216,217,217,218,218,218,218,218,219,220,221,220,221,221,221,221,221,220,220,220,221,221,221,220,219,218,218,218,218,217,217,218,218,217,216,217,217,215,215,214,214,213,212,212,212,213,212,212,211,211,211,209,209,209,208,208,208,207,206,205,204,205,205,202,202,204,204,202,202,203,201,202,200,201,199,199,201,200,199,200,200,200,201,200,200,201,200,204,198,199,198,200,200,193,193,196,196,195,196,197,197,197,199,199,200,201,202,202,203,205,205,206,208,208,208,209,210,211,211,211,212,213,213,214,215,215,215,215,215,215,216,217,218,218,217,218,217,217,218,220,220,219,220,220,221,221,221,221,220,220,221,221,221,221,220,219,219,220,220,219,218,219,219,218,217,217,217,216,216,216,215,214,214,214,214,214,213,212,212,212,212,210,211,210,209,209,209,208,208,207,206,206,205,204,203,204,204,203,204,204,202,204,201,202,199,200,202,200,201,202,200,201,202,200,200,199,200,203,200,200,201,203,203,193,193,196,197,195,196,197,196,196,199,199,201,202,203,203,204,205,206,207,208,209,209,209,210,212,212,213,213,213,214,214,214,215,215,215,215,215,216,217,218,219,218,218,218,218,219,220,220,219,220,220,220,221,221,221,221,221,221,221,222,221,220,220,220,221,221,219,218,219,219,218,217,217,217,217,217,216,215,214,214,214,215,215,214,212,211,212,212,211,212,211,209,208,208,208,208,208,208,206,206,206,205,204,205,206,204,205,202,204,202,204,201,201,202,199,201,203,199,201,202,198,201,199,203,202,201,196,201,203,203,197,197,195,196,196,196,198,200,199,200,202,203,202,203,205,206,206,206,209,210,209,210,210,210,211,210,211,213,214,214,214,215,215,217,217,217,216,216,217,218,218,217,217,218,218,219,219,220,220,219,220,220,220,221,222,222,221,221,221,221,221,220,220,220,220,220,220,220,220,220,219,218,218,218,218,217,216,216,216,215,214,214,214,214,214,213,212,212,213,212,212,211,212,212,212,207,211,205,211,207,204,209,207,204,206,204,206,202,203,201,204,202,201,202,202,202,202,202,202,202,202,203,202,203,203,202,200,201,204,204,196,196,195,196,197,197,198,200,200,201,202,203,203,204,205,205,205,207,209,209,210,211,211,211,213,211,212,214,215,215,215,216,216,216,217,217,216,216,217,218,219,218,218,219,219,220,220,220,220,220,220,221,221,222,222,222,221,221,221,221,221,221,221,221,221,221,221,221,220,220,219,218,217,218,218,217,216,216,215,215,214,215,214,213,214,214,213,212,212,211,213,212,209,210,209,215,208,212,203,206,208,201,184,206,204,203,206,203,206,202,203,201,202,202,202,203,203,202,202,202,202,202,201,202,202,201,199,200,203,203,195,195,195,196,198,198,199,201,201,200,202,203,204,205,207,207,207,208,209,209,210,212,212,211,214,213,213,214,215,215,216,217,217,217,217,218,217,217,218,219,219,219,219,220,220,220,221,221,221,221,221,221,221,222,222,222,221,221,221,221,221,221,221,221,221,222,221,221,220,220,219,218,217,218,218,218,216,215,215,214,214,215,213,212,213,214,214,212,211,210,212,211,212,212,212,210,212,203,198,207,205,202,165,192,204,208,200,205,204,204,205,203,204,202,203,203,203,203,202,202,202,202,202,202,202,200,199,200,202,202,195,195,195,197,199,199,200,202,202,201,202,202,203,205,207,207,207,209,210,210,211,212,212,211,214,213,214,214,215,215,216,217,217,217,218,218,218,218,219,220,220,220,220,220,221,221,221,221,221,221,221,221,221,221,222,221,221,221,221,221,221,221,221,221,221,221,221,221,220,220,219,218,218,218,218,218,216,215,215,214,214,214,212,212,213,214,214,213,211,213,210,210,213,211,208,206,210,186,210,200,208,198,183,174,191,188,207,201,205,205,208,202,204,202,203,204,204,203,202,202,203,203,202,202,202,200,199,200,201,201,196,196,196,198,200,200,201,202,202,203,203,202,203,204,205,206,206,208,210,210,211,212,212,212,213,214,214,214,215,215,216,217,217,218,219,220,219,219,220,221,221,221,221,221,221,221,221,221,221,221,221,221,221,220,221,220,220,220,220,220,221,221,220,220,220,220,220,220,220,219,219,218,218,217,218,218,216,215,214,214,214,212,212,212,213,213,213,212,212,211,211,210,210,210,206,214,211,206,148,183,191,176,186,175,186,154,204,181,200,203,208,201,204,203,204,204,204,203,202,202,203,202,202,202,201,200,199,199,200,200,198,198,198,200,201,200,201,202,202,204,203,202,203,205,206,208,209,206,210,211,211,212,213,213,214,214,214,214,215,216,217,218,218,219,220,220,220,220,221,221,221,221,221,221,221,221,221,221,221,220,221,221,220,220,220,220,220,220,220,220,220,220,220,220,220,220,220,220,219,218,218,217,217,217,218,217,216,214,214,213,213,212,212,212,212,212,211,211,211,208,213,212,211,207,209,187,211,214,165,171,173,165,170,169,167,178,179,173,189,202,207,203,206,204,204,204,203,202,202,203,203,203,203,202,201,200,199,200,200,200,199,199,199,201,202,200,201,202,202,204,203,203,205,206,207,209,212,205,212,214,211,212,215,215,214,214,214,214,215,217,218,218,218,218,220,220,220,220,220,221,221,221,221,221,221,221,221,221,221,221,221,221,220,220,220,220,220,220,220,220,220,220,220,220,219,219,219,219,218,218,217,217,217,217,217,216,215,214,214,213,212,211,211,210,210,210,210,209,210,209,212,210,210,196,191,158,195,200,172,173,169,173,157,155,159,205,169,192,194,204,205,204,204,205,204,203,202,202,202,203,203,203,203,202,201,200,200,200,200,200,198,198,198,201,202,200,201,203,203,205,204,205,206,206,205,207,209,205,213,215,212,212,215,215,213,213,213,214,215,217,217,217,217,218,219,220,220,220,220,220,220,221,221,221,221,221,221,221,221,221,222,222,221,220,220,220,220,220,220,221,221,220,220,220,219,218,218,218,217,217,217,217,217,217,216,215,214,213,213,212,211,211,209,209,209,209,209,209,210,209,207,208,206,188,167,179,185,194,182,172,171,165,168,154,173,166,172,204,207,202,202,204,205,205,204,203,202,202,202,203,203,202,202,201,200,199,199,199,199,199,200,200,196,203,202,202,201,204,204,206,205,204,208,209,204,213,204,105,210,211,211,213,215,215,214,214,215,212,215,219,214,219,218,220,220,220,219,220,220,220,220,220,221,221,221,221,221,221,221,221,222,222,222,220,220,220,221,217,221,218,223,220,219,220,219,219,218,218,218,217,216,216,218,216,215,215,215,215,213,212,212,212,207,209,208,212,209,208,208,212,210,202,189,198,186,173,173,168,197,167,166,169,155,157,154,172,178,180,203,202,204,201,205,207,204,205,202,202,203,202,202,201,202,202,203,203,199,197,199,199,199,199,195,202,202,202,202,204,204,205,204,208,206,203,209,210,164,182,197,184,216,212,214,212,214,217,214,216,218,215,219,216,218,219,220,220,220,220,221,221,221,221,221,221,221,221,221,221,221,221,222,222,222,221,220,220,221,222,221,219,218,217,220,224,216,219,218,217,218,217,216,217,218,216,215,215,215,215,214,212,212,210,211,212,210,207,207,211,209,206,204,210,187,176,183,174,179,173,157,176,170,165,163,153,155,204,166,203,205,200,203,205,204,203,205,203,204,203,204,203,203,203,203,203,203,203,200,197,199,199,198,198,195,201,202,202,202,205,205,207,206,204,206,209,209,207,174,129,141,175,175,211,215,213,217,212,217,219,214,221,218,218,218,217,219,220,220,220,220,221,221,221,221,221,221,221,221,221,222,221,222,222,222,222,221,221,220,219,220,221,217,223,221,219,223,220,219,218,217,217,216,216,217,215,215,215,215,215,215,213,212,211,213,206,209,213,210,207,206,215,199,209,179,178,178,169,179,169,159,167,166,166,158,161,151,203,190,197,205,203,203,202,205,206,208,201,205,202,203,204,204,203,203,203,204,205,202,200,202,202,198,198,194,201,201,202,203,205,205,206,204,209,205,205,204,197,121,115,126,176,174,218,210,214,213,219,212,212,218,215,220,217,215,216,218,220,220,220,220,220,220,221,221,221,221,222,222,223,223,223,223,223,224,224,223,221,220,221,217,223,222,219,221,218,218,220,219,218,217,217,216,215,215,215,215,215,215,215,215,214,212,211,212,209,211,211,211,210,212,209,182,172,163,171,164,175,161,152,160,164,166,170,161,157,154,199,199,203,207,202,201,203,204,200,203,195,206,204,204,203,201,203,203,202,203,205,204,202,203,203,198,198,194,201,201,202,202,205,204,204,207,207,207,199,210,131,120,107,117,97,209,212,208,208,207,213,213,206,220,213,218,221,213,217,219,220,220,220,220,220,220,221,221,221,221,222,222,223,223,223,223,224,224,224,223,221,219,219,217,216,219,218,221,220,223,218,218,218,218,217,217,216,215,215,215,215,215,215,215,214,213,212,209,215,213,209,212,209,205,208,207,199,170,166,163,159,161,151,150,166,172,166,151,148,157,200,193,196,187,198,201,203,200,204,203,193,205,203,202,203,203,203,203,202,202,204,203,201,202,202,200,200,195,202,202,203,203,205,204,206,207,203,203,207,207,148,141,124,126,122,208,149,157,213,147,152,206,111,217,219,212,209,216,217,219,220,220,220,220,220,220,221,221,221,221,221,221,221,221,222,222,222,222,222,221,219,218,217,172,83,209,225,212,223,214,217,217,218,218,218,218,218,217,217,218,218,217,217,217,216,214,214,214,214,209,214,211,210,215,211,213,208,204,178,202,166,154,158,153,161,168,164,139,148,150,191,195,200,165,195,199,198,200,199,199,194,202,201,202,203,204,202,203,202,202,203,203,202,203,203,200,200,195,201,202,203,203,205,204,207,204,208,207,199,210,203,209,106,203,129,180,118,147,205,157,169,200,139,216,215,220,194,215,216,218,219,219,219,220,220,219,220,220,221,221,221,220,220,220,220,220,220,221,221,220,219,218,214,85,30,138,195,224,218,221,218,219,219,218,218,219,219,218,219,220,220,218,218,219,218,216,215,218,215,209,214,209,217,207,207,213,208,202,206,191,190,156,152,153,162,163,163,148,144,144,186,168,195,164,198,199,198,175,170,182,193,201,202,203,201,199,200,202,201,201,203,203,203,205,205,198,198,194,200,200,202,202,204,203,203,206,208,207,205,206,203,212,174,200,123,121,124,133,204,199,191,98,115,191,197,209,199,212,215,216,217,217,218,219,219,219,220,220,221,221,221,221,221,220,220,221,221,222,222,221,221,220,94,109,40,53,84,162,214,215,220,221,220,219,218,219,220,219,220,221,220,218,217,219,218,216,218,211,216,216,214,215,212,134,215,209,204,193,180,186,195,172,154,160,161,166,150,141,143,143,133,141,160,189,184,164,186,165,166,182,198,197,196,200,201,201,199,201,200,199,200,201,201,202,202,197,197,197,201,201,200,204,205,201,204,208,205,206,204,207,192,206,181,161,112,128,115,129,114,142,158,135,119,128,158,43,129,215,214,222,217,215,220,219,218,222,220,220,220,220,221,222,222,221,223,218,222,221,221,221,222,212,129,37,25,104,167,143,156,194,216,224,218,222,219,218,221,221,220,221,217,218,222,217,218,218,218,215,216,213,213,216,211,163,212,216,170,180,168,185,151,154,151,152,157,165,156,141,148,119,123,134,108,152,151,157,156,161,174,198,162,198,197,200,200,199,201,201,200,199,199,198,200,203,203,202,202,193,199,205,198,199,205,204,202,206,206,209,204,123,174,176,178,156,90,124,93,128,122,148,171,148,142,142,137,138,140,218,215,220,220,221,222,221,225,219,220,221,222,221,221,220,220,219,217,221,220,223,223,223,225,210,80,60,101,172,123,133,191,153,167,218,211,218,221,224,219,220,219,220,222,219,216,216,218,216,217,216,214,219,216,213,207,167,201,207,170,164,142,134,140,160,146,155,160,167,152,144,148,146,142,126,117,151,148,155,152,162,182,160,193,196,193,198,199,200,197,198,200,199,202,198,198,200,200,192,192,198,199,198,199,201,202,201,205,199,205,206,205,163,133,146,174,159,86,113,96,105,110,152,170,165,151,139,148,161,156,187,218,217,222,220,222,217,215,222,221,221,221,220,219,221,223,225,223,225,223,221,225,229,205,142,34,64,144,174,201,165,91,181,168,176,206,224,221,219,221,217,221,222,216,217,222,213,219,213,209,216,211,206,211,208,205,161,187,181,164,156,158,135,151,153,140,148,160,156,160,143,146,154,159,144,145,144,148,151,148,163,159,183,191,189,192,194,199,191,197,192,197,194,195,197,198,201,201,195,195,198,196,199,204,198,196,202,196,202,202,207,209,206,198,148,152,154,57,92,92,99,106,136,160,167,157,153,148,154,156,166,221,218,224,219,213,219,222,220,220,220,222,223,223,222,221,221,223,222,221,222,220,216,146,57,57,93,178,177,180,215,208,160,183,186,184,189,220,222,215,220,217,219,217,213,209,207,211,219,216,209,211,207,202,188,178,86,174,176,166,165,164,140,145,144,136,152,163,158,158,141,144,156,148,142,143,151,144,143,147,146,147,158,162,164,195,201,194,195,195,195,198,199,196,200,199,197,197,199,199,193,193,202,202,202,204,197,200,198,137,86,198,211,193,153,155,104,59,64,85,99,120,132,140,157,167,162,85,142,166,182,220,223,216,219,218,218,222,221,225,223,222,222,223,222,222,223,222,222,221,220,217,197,39,59,72,169,179,230,191,208,104,163,177,190,192,191,188,183,210,214,215,213,216,210,174,155,165,172,145,144,146,144,149,133,96,23,163,177,171,161,163,143,178,143,146,152,156,148,161,143,155,150,150,144,143,137,126,152,118,106,128,184,197,192,195,200,198,194,198,203,197,200,195,200,203,198,198,192,192,193,195,199,200,205,198,169,162,160,104,103,201,178,122,146,159,161,165,93,117,107,107,122,116,127,154,160,137,40,104,188,216,218,222,221,223,223,221,226,221,219,218,219,219,218,218,220,216,206,208,197,204,157,120,65,139,176,203,216,231,164,53,152,121,187,194,193,195,191,187,121,137,123,121,112,155,164,173,170,163,169,162,172,177,169,109,70,54,171,168,157,166,160,163,136,142,153,140,157,146,144,152,152,142,140,136,114,86,116,136,104,131,168,164,168,199,200,200,200,203,172,198,192,168,199,198,196,196,195,195,194,194,200,201,199,180,137,144,150,107,113,98,93,88,140,131,160,175,157,95,73,99,102,106,89,132,141,60,93,142,132,220,221,225,219,223,221,226,216,210,201,188,177,170,170,175,182,182,181,193,186,173,117,49,137,177,190,218,215,227,212,216,216,205,98,185,195,198,193,186,170,156,94,110,116,149,163,167,174,172,167,171,160,170,168,47,82,59,124,176,157,171,170,161,142,151,146,126,153,154,149,150,146,139,129,132,119,115,114,134,119,154,187,168,197,197,201,199,203,189,195,187,188,196,190,191,200,200,193,193,192,196,197,192,206,191,125,137,143,109,109,83,94,76,144,124,159,169,155,125,41,27,51,44,105,127,129,97,116,152,116,208,218,171,179,217,164,166,173,175,178,182,186,187,185,187,191,184,193,192,153,118,28,66,173,176,202,205,225,214,227,216,213,203,209,181,189,192,194,190,190,179,154,101,112,113,141,160,172,169,173,161,164,164,146,80,169,141,47,166,167,173,167,164,158,158,143,117,150,154,148,142,145,143,133,135,125,118,112,129,148,155,203,184,202,200,200,198,196,187,197,184,179,199,179,178,194,194,191,191,195,197,200,194,180,133,121,137,142,135,95,69,97,74,143,129,152,152,119,106,84,13,1,32,23,66,80,80,118,158,173,215,191,146,159,203,184,183,178,180,181,184,192,186,186,187,189,192,189,180,77,34,56,57,181,193,229,212,219,222,228,225,209,223,171,109,182,190,193,186,189,194,181,150,67,105,113,153,169,168,174,165,163,160,46,87,88,196,45,162,171,171,170,166,163,155,153,107,146,150,144,134,133,141,146,123,125,110,121,127,151,149,177,201,197,202,198,204,193,187,198,182,183,184,182,170,177,177,197,197,195,196,197,187,134,138,144,147,151,146,106,94,87,75,88,89,130,141,87,95,66,57,55,88,62,83,62,47,64,146,185,160,151,140,163,185,195,193,190,192,190,185,190,190,186,187,191,190,183,122,109,58,143,182,192,202,213,224,206,224,224,223,215,216,213,192,68,187,190,191,190,192,183,175,117,91,140,136,165,172,164,161,158,155,95,81,82,144,87,76,172,171,174,167,163,166,166,142,138,113,149,121,133,142,154,117,126,127,125,115,143,149,163,194,183,202,201,189,198,187,189,189,184,183,181,174,193,193,193,193,192,198,195,177,116,120,144,145,165,153,116,103,102,88,87,91,209,177,71,80,68,64,65,87,98,91,96,35,35,117,158,167,148,154,163,185,188,197,192,191,189,192,195,192,186,188,190,185,164,133,42,54,160,187,187,217,221,226,220,227,226,226,222,206,220,214,222,139,188,183,185,187,179,163,145,86,136,146,165,163,170,165,163,115,99,87,87,39,173,40,162,174,176,164,161,162,144,138,121,130,143,143,134,137,130,140,136,129,124,128,117,129,146,177,166,183,192,184,190,185,189,184,185,186,180,192,198,198,199,199,199,195,179,176,122,130,126,186,172,159,150,96,98,97,92,92,74,75,47,64,66,75,69,77,82,111,114,116,147,148,149,149,152,144,153,89,187,196,188,190,186,189,187,191,191,189,188,182,74,91,52,119,180,189,212,213,220,212,231,223,227,228,226,211,213,216,149,155,155,179,179,179,167,159,185,152,69,133,181,169,163,164,154,98,85,120,110,91,69,66,128,167,170,157,141,122,122,145,120,135,143,143,138,135,144,140,149,141,128,133,133,120,134,157,139,152,190,188,186,190,187,188,184,187,197,200,197,197,197,197,193,199,188,195,193,195,156,135,165,161,134,103,104,106,84,71,84,41,79,73,60,65,63,58,61,86,91,140,158,166,167,137,153,138,66,83,190,189,193,192,189,191,185,190,189,183,182,159,106,48,56,168,181,188,226,225,218,224,231,227,227,223,225,222,204,211,219,148,111,174,190,198,183,170,178,164,74,140,180,168,166,163,53,118,85,133,136,81,39,194,48,169,148,133,152,115,75,114,143,138,141,141,140,143,139,146,145,142,133,135,139,133,141,128,136,143,197,188,186,188,187,184,183,184,201,197,188,188,199,199,195,199,199,201,205,194,197,126,133,147,119,106,102,101,78,74,77,46,83,76,57,66,58,60,48,59,111,115,134,156,161,126,44,148,168,179,198,186,192,193,184,189,189,183,188,188,168,115,54,57,119,178,177,214,217,224,212,226,223,228,225,227,226,224,207,225,87,84,128,83,183,178,179,178,160,149,107,75,172,162,164,146,101,87,102,108,138,117,87,81,24,128,133,122,172,102,118,139,143,130,135,152,139,139,145,141,144,140,131,138,132,123,125,130,129,187,191,182,184,187,187,172,185,185,195,190,179,179,198,198,194,198,200,199,202,206,139,170,124,123,109,102,105,93,81,77,71,68,114,96,54,50,51,40,44,36,87,96,115,124,151,113,173,154,145,191,200,144,156,192,195,187,187,178,184,179,124,45,21,20,166,169,210,231,203,227,224,224,227,226,225,229,222,223,226,204,213,195,56,93,74,92,167,171,171,116,113,74,149,163,159,137,137,71,105,127,138,113,99,43,29,76,103,120,164,121,126,134,136,129,136,136,133,139,129,135,132,139,119,128,134,109,119,123,124,124,193,203,180,191,185,177,184,184,196,178,182,182,194,194,199,196,198,202,202,190,119,140,114,101,99,106,102,87,85,74,82,36,156,140,51,33,61,36,30,43,94,93,85,89,126,144,144,148,157,195,176,162,152,132,191,189,190,192,189,171,111,140,70,112,180,186,196,224,230,224,226,224,229,225,231,231,223,224,225,221,215,210,128,65,19,52,64,123,116,146,115,117,136,142,145,76,90,86,123,124,141,122,106,89,25,35,123,69,152,123,126,145,134,130,124,125,135,128,137,126,141,140,135,126,133,112,114,104,121,151,121,197,167,182,189,178,184,179,181,175,181,181,197,197,195,201,198,201,125,118,111,105,125,73,96,98,108,83,82,74,41,18,85,126,50,48,95,74,44,81,98,110,78,32,71,137,139,130,165,160,182,181,194,171,182,198,200,204,206,75,30,92,194,195,193,204,188,227,232,232,229,225,228,231,231,230,230,228,222,226,222,216,149,165,50,24,24,71,75,50,128,134,111,136,156,113,84,101,135,145,159,125,144,107,44,10,89,134,83,138,158,139,150,146,133,116,126,137,126,77,145,144,130,130,134,115,111,122,133,136,134,153,179,187,185,185,184,180,178,170,183,183,196,196,199,195,205,194,123,111,116,132,102,50,76,107,106,94,85,78,16,45,146,20,92,65,128,126,96,85,84,122,107,165,25,135,134,120,111,131,147,187,194,151,161,195,192,195,207,65,152,183,150,184,202,233,182,200,222,232,233,223,223,227,228,226,233,227,221,225,224,212,147,146,124,112,43,43,41,62,98,33,132,149,99,82,86,115,142,152,160,121,150,136,81,21,29,158,102,92,113,110,148,162,127,121,118,126,125,125,117,143,137,131,134,125,108,137,137,136,119,157,173,179,180,187,187,182,185,179,181,181,198,198,196,203,197,203,124,108,118,96,87,73,57,85,105,99,84,73,65,60,108,145,87,111,157,104,82,74,61,109,113,133,71,131,112,76,37,44,125,152,179,105,198,196,184,192,213,191,191,205,207,181,225,213,237,225,221,229,231,227,227,223,225,228,228,231,225,221,224,204,132,128,124,120,127,125,89,76,44,42,59,57,72,28,103,142,143,143,152,121,131,145,90,32,65,120,150,68,102,112,111,156,131,85,117,125,144,136,68,141,94,139,131,109,123,135,198,192,172,183,185,188,185,187,183,177,185,186,186,186,198,198,201,67,79,171,158,119,146,105,107,78,65,56,74,90,87,71,75,51,60,141,58,69,37,22,47,16,80,79,96,108,130,126,107,93,190,137,81,88,189,164,153,189,192,189,204,204,195,209,198,194,229,213,229,225,221,225,232,226,227,229,224,225,231,227,227,224,217,219,170,130,115,123,123,149,150,140,66,54,87,21,63,34,137,146,134,131,136,113,119,111,89,59,54,32,118,100,113,104,122,143,132,94,107,99,126,136,101,79,132,132,133,90,116,129,147,130,177,189,189,193,188,190,187,182,184,184,184,184,198,198,196,94,84,139,134,152,121,110,114,101,86,59,83,94,67,62,82,40,61,121,52,40,183,99,93,133,77,105,91,84,125,142,145,146,116,94,106,127,152,155,198,206,209,207,207,210,195,214,203,208,222,228,214,229,227,225,234,227,225,226,230,233,229,230,228,220,222,221,192,139,103,121,117,122,119,138,117,108,128,49,20,57,141,142,111,124,126,98,102,136,86,78,66,3,53,107,116,138,137,138,96,109,108,107,115,123,125,76,135,141,110,77,98,127,126,88,186,193,188,188,190,191,188,189,186,182,183,183,189,189,153,48,196,185,157,118,95,85,101,88,74,46,90,71,74,57,71,52,46,113,151,22,132,130,102,169,76,117,70,70,147,149,171,115,93,72,145,80,80,187,202,199,189,186,180,175,159,214,97,223,196,225,223,229,226,228,233,217,227,232,234,227,226,228,224,225,221,223,193,133,97,110,113,117,114,144,107,106,127,101,47,75,140,105,93,93,123,93,79,110,117,68,63,6,17,140,95,74,74,136,91,107,114,110,110,121,105,131,138,142,82,72,56,125,132,159,194,189,198,189,194,191,184,188,188,186,185,185,197,197,199,119,119,202,175,101,85,74,66,54,114,59,72,46,55,45,38,45,46,40,219,29,111,83,92,154,106,74,75,127,73,84,110,53,169,128,170,190,170,202,211,159,85,45,43,53,51,94,129,218,178,231,234,230,225,221,231,176,169,184,223,222,228,228,224,223,225,219,177,139,93,110,109,115,108,129,110,105,127,99,51,95,130,99,90,90,114,81,71,67,107,73,63,17,74,166,54,136,27,97,71,101,108,113,89,110,96,130,126,106,70,66,62,123,161,199,171,187,187,189,192,193,189,191,188,188,183,183,192,192,194,174,39,207,134,72,86,56,60,63,76,69,64,51,40,11,17,30,43,40,180,139,110,83,57,102,40,69,56,22,67,112,191,140,58,40,52,61,57,57,92,68,53,70,131,63,58,97,100,218,219,231,230,226,227,223,191,145,176,168,214,227,229,228,226,222,221,222,193,139,137,112,106,112,108,131,106,99,130,98,58,81,119,104,79,88,93,37,43,82,155,189,130,158,170,153,152,124,35,88,85,81,128,110,104,94,105,113,130,100,61,86,67,89,134,102,128,179,189,192,188,192,192,191,185,188,184,184,171,171,197,126,51,200,104,78,98,74,52,76,80,79,62,46,21,9,16,40,46,44,93,129,114,89,51,37,81,84,57,49,60,20,26,67,85,66,76,92,77,78,103,133,134,131,158,123,145,147,137,215,221,229,235,224,228,204,169,92,72,150,186,226,228,230,227,223,222,220,210,117,141,138,127,112,113,123,100,103,131,99,53,71,104,78,98,128,77,63,116,143,179,189,158,147,156,178,164,48,95,99,75,71,107,80,89,83,87,97,119,63,77,79,72,66,91,83,131,170,186,191,194,186,193,188,185,186,186,186,106,106,193,184,204,197,161,117,188,45,67,72,81,76,58,44,20,40,33,166,44,44,67,82,126,81,60,21,107,73,67,55,41,37,44,55,135,147,133,151,131,134,133,158,167,152,145,112,155,177,161,211,232,231,231,231,207,196,97,79,94,114,170,207,227,228,222,224,223,222,212,112,135,150,146,134,131,116,89,89,140,99,54,74,97,94,107,116,145,115,135,138,172,195,155,111,165,174,96,157,68,89,47,40,70,61,81,68,86,81,98,81,88,74,60,71,101,102,128,172,177,191,191,190,189,188,184,184,184,184,154,154,179,198,198,190,199,197,162,58,72,77,70,60,42,41,19,57,59,113,47,47,50,68,157,77,72,56,74,24,14,10,25,46,61,79,94,111,160,167,132,167,133,131,142,118,131,148,155,154,166,210,226,226,225,223,194,166,72,55,128,127,206,182,219,227,217,227,222,221,215,107,131,127,106,120,112,100,104,106,109,108,62,74,49,81,98,99,126,128,128,146,177,183,161,156,158,127,56,69,136,46,51,21,72,60,72,68,66,75,73,77,76,84,57,93,113,126,129,162,176,184,183,188,183,184,184,180,183,183,131,131,133,178,164,197,196,86,76,68,63,79,72,58,18,54,32,118,95,67,43,41,52,68,161,80,95,82,68,23,11,13,30,80,137,127,106,116,91,73,97,137,157,162,168,160,163,171,160,160,169,213,227,230,228,223,188,111,52,74,204,183,91,154,220,222,223,221,223,222,213,121,133,116,112,120,126,114,105,111,106,105,62,52,49,90,98,104,104,127,143,154,185,169,159,156,161,50,55,121,118,45,41,42,51,72,70,73,66,68,75,86,77,58,81,109,92,154,135,161,174,178,178,186,179,181,186,177,182,182,142,142,133,178,158,183,121,86,74,81,64,72,74,70,53,46,153,132,76,56,58,31,47,57,178,76,106,79,30,17,42,69,72,76,90,90,95,109,136,151,147,163,163,167,166,163,166,160,151,155,168,222,229,221,229,225,116,48,46,216,224,224,121,190,203,220,223,224,222,221,221,129,141,105,117,128,119,120,113,110,111,93,53,49,46,100,106,110,127,132,130,171,185,166,156,153,153,78,123,123,120,107,56,54,20,68,88,84,65,66,70,84,94,209,107,106,189,192,122,166,166,178,178,187,175,183,186,177,178,178,117,117,134,162,152,124,113,73,76,79,60,50,59,68,54,90,131,105,35,90,110,19,36,48,102,68,60,62,24,77,66,66,68,70,76,80,113,107,134,152,147,159,161,154,151,154,149,145,147,154,158,227,226,230,227,223,177,38,109,232,223,219,216,142,172,220,222,226,221,219,221,126,136,123,104,111,118,116,127,119,97,98,57,46,87,98,114,113,124,140,142,170,167,149,149,144,86,83,110,102,111,127,36,68,40,59,82,66,71,45,88,71,83,193,174,197,190,182,172,153,163,172,172,182,167,185,183,181,175,175,124,124,114,144,126,112,101,80,69,55,45,44,59,55,46,100,119,108,32,128,82,152,75,37,88,54,77,55,26,80,82,70,72,85,89,90,121,111,141,142,126,139,155,144,145,151,149,154,150,146,156,226,227,226,224,226,155,50,34,64,121,135,89,209,214,219,228,218,224,221,209,126,123,106,87,54,95,129,107,93,111,111,59,30,99,96,86,113,137,143,146,156,147,151,150,124,70,79,99,112,89,149,115,61,62,30,71,70,65,46,84,68,85,83,102,195,165,177,166,162,164,158,165,167,160,181,183,184,174,174,128,128,128,140,116,106,98,75,68,83,40,60,115,51,56,144,129,43,15,135,133,133,135,99,49,64,31,54,134,83,76,79,71,82,95,100,122,118,141,138,135,144,148,150,153,150,154,155,147,137,131,229,227,226,226,224,222,143,154,159,143,141,61,222,217,224,218,226,222,219,217,114,125,102,37,48,49,121,112,115,101,112,31,63,99,40,84,120,138,144,154,153,151,145,156,40,75,71,91,91,118,124,129,14,34,34,76,68,62,52,73,77,67,135,101,186,149,172,171,153,152,150,163,154,161,175,186,183,174,174,134,134,169,144,150,100,89,61,66,119,45,86,63,53,61,104,124,104,61,15,110,99,32,61,61,68,47,59,49,74,77,67,61,57,75,100,116,130,144,137,137,146,145,153,134,132,124,134,137,169,144,223,226,226,226,223,219,166,152,146,149,129,59,216,219,223,224,224,222,221,214,122,120,46,72,64,42,133,91,59,49,92,38,98,110,92,109,143,142,150,157,152,154,168,90,47,98,110,96,82,116,128,125,102,5,39,38,78,47,74,101,90,85,84,111,113,195,175,157,150,151,162,157,157,166,178,184,183,173,173,127,127,121,149,116,111,91,85,56,60,78,100,54,57,54,107,106,106,145,110,58,31,27,80,91,68,40,7,13,94,85,80,95,90,130,134,123,117,57,111,43,162,118,192,202,199,202,201,208,205,210,220,227,224,227,228,224,150,157,148,141,99,94,210,221,222,223,223,222,221,214,119,122,45,97,110,23,197,57,53,40,37,83,103,96,100,121,137,157,165,156,159,169,166,74,108,131,136,111,84,108,129,111,136,18,26,30,94,43,91,101,91,82,86,97,153,201,148,161,145,152,150,165,154,161,186,185,180,166,166,121,121,133,137,55,162,77,98,85,95,87,78,53,38,79,110,92,105,76,71,28,39,25,30,57,35,10,46,101,126,112,78,113,182,157,181,166,186,208,194,201,205,206,205,205,209,208,203,206,208,209,219,224,232,221,225,212,153,154,154,142,57,106,191,223,221,221,222,223,221,216,116,126,65,98,92,24,58,33,40,44,26,101,106,56,82,131,153,167,167,147,168,174,24,17,80,123,139,100,78,129,136,130,138,70,58,58,48,85,100,92,86,81,88,95,168,104,126,151,152,147,149,157,151,159,177,183,171,168,168,124,124,131,142,33,134,131,84,100,97,113,76,60,17,58,82,66,70,33,16,22,20,33,24,74,53,126,142,113,128,133,152,163,202,201,194,203,198,202,201,205,206,199,207,205,207,205,205,212,215,206,218,227,223,229,225,144,154,151,159,138,85,101,157,220,222,221,221,223,220,215,113,128,85,146,130,11,47,43,65,46,61,77,80,24,76,155,155,112,156,130,61,34,93,44,119,115,114,123,102,124,121,125,132,123,67,53,53,59,169,88,98,112,145,109,169,198,150,153,153,148,148,148,154,157,181,172,170,161,161,125,125,138,139,140,142,144,197,165,149,93,64,34,25,29,52,29,37,68,13,14,19,29,25,142,144,133,133,151,145,167,163,168,200,198,198,192,201,196,205,202,203,204,207,204,202,209,212,206,211,95,220,224,225,227,231,159,121,87,46,67,63,90,159,218,220,220,221,223,222,220,119,136,109,173,171,151,66,81,35,83,32,25,27,25,28,38,50,59,57,56,30,29,39,46,123,122,133,121,109,142,133,129,133,118,91,40,29,96,97,104,104,137,134,98,147,121,118,154,141,147,150,152,154,151,176,171,164,162,162,123,123,140,149,146,144,135,103,91,63,65,55,59,29,14,11,15,19,9,16,10,10,17,77,170,150,145,150,102,62,132,155,194,203,195,194,191,201,199,200,203,203,201,202,212,202,206,203,211,206,73,204,229,227,223,227,206,136,19,27,33,26,32,161,224,223,222,220,219,217,212,113,124,62,93,80,161,96,102,46,54,70,41,44,39,42,28,101,61,137,93,45,42,41,61,123,136,143,137,109,144,137,136,138,116,81,45,23,102,130,136,134,102,77,145,96,170,136,206,190,142,147,150,152,161,173,162,164,167,167,122,122,140,142,142,148,143,58,95,60,70,40,96,14,12,5,79,64,14,11,9,6,175,155,159,95,100,102,53,76,168,189,199,196,193,195,198,194,197,206,195,201,204,209,204,197,194,201,189,38,58,195,229,222,214,221,226,135,20,201,27,32,44,171,208,220,220,221,221,222,218,126,130,51,97,52,153,108,102,54,79,99,100,99,65,50,56,108,59,144,114,94,72,58,93,117,145,148,138,109,145,142,128,148,100,84,51,33,116,153,145,145,123,111,180,130,180,200,159,146,141,146,147,145,168,175,158,163,174,174,132,132,148,148,140,150,67,62,105,47,203,69,216,26,50,130,136,145,139,146,156,38,188,186,109,105,129,87,56,149,195,200,195,189,192,193,192,195,198,184,196,204,201,202,200,181,200,185,103,89,63,171,227,223,201,221,222,138,20,162,39,46,29,170,184,221,222,222,220,220,215,124,123,64,49,44,137,113,99,48,73,103,59,101,78,74,91,107,53,140,122,78,69,75,124,125,140,161,127,117,147,145,145,140,96,98,50,67,124,167,149,159,147,156,153,152,159,170,164,158,146,141,142,155,179,149,161,52,85,85,133,133,161,114,138,144,53,42,65,154,12,135,184,178,145,149,139,135,150,163,152,183,199,101,54,66,73,55,74,192,191,191,186,187,189,193,195,190,193,206,154,199,185,201,188,184,188,112,79,92,52,175,224,223,191,225,208,153,16,87,31,49,30,173,165,219,223,220,220,220,216,125,126,67,63,48,150,114,106,52,70,102,84,94,84,84,82,134,61,143,107,120,123,158,165,131,139,162,143,120,147,129,129,149,113,101,58,89,136,146,153,159,152,150,153,167,168,171,173,153,153,148,142,159,170,129,151,78,82,82,145,145,151,82,155,83,43,44,145,161,134,161,187,152,183,161,157,133,124,161,190,198,155,46,50,49,52,70,170,188,185,186,183,184,185,189,193,195,173,56,155,171,74,116,218,176,156,111,83,93,63,192,227,226,199,219,209,172,27,45,24,31,41,171,168,221,221,221,221,221,215,127,124,82,70,54,134,118,118,60,88,116,41,132,72,82,98,141,63,137,109,125,172,169,162,121,146,141,119,124,121,138,127,147,151,119,58,107,142,148,144,165,158,157,153,161,179,178,173,166,148,152,157,171,158,136,137,108,133,133,134,134,92,75,152,114,143,119,156,160,150,171,128,177,174,167,161,158,154,180,196,173,53,49,52,84,137,176,191,191,174,175,173,176,175,182,34,79,86,86,72,87,95,62,74,140,146,68,77,69,64,197,221,226,198,220,210,186,45,118,137,134,142,180,173,221,221,222,220,220,215,131,126,97,90,49,133,129,124,69,80,107,37,130,139,117,123,156,64,137,101,127,198,203,194,124,149,141,127,126,131,118,122,132,150,108,65,127,184,155,152,173,166,165,150,157,179,177,177,170,131,137,172,162,145,139,127,124,122,122,96,96,75,74,77,135,82,145,147,135,117,172,188,184,172,175,168,167,168,188,176,47,47,43,66,107,188,132,141,170,165,173,153,80,40,45,107,101,102,105,107,116,113,100,90,129,142,66,68,58,46,166,212,224,172,223,207,210,180,133,184,186,172,182,176,204,220,222,220,219,214,128,126,112,70,53,124,133,127,57,75,92,44,108,144,138,122,153,91,96,112,177,206,205,202,97,150,135,138,126,128,128,129,129,151,125,72,57,207,191,200,160,182,179,162,167,176,162,138,163,130,124,165,134,137,121,132,135,120,120,74,74,78,72,65,87,92,162,147,109,142,194,186,187,181,166,159,168,181,168,88,77,79,81,89,76,38,50,40,45,58,72,66,97,105,104,124,124,122,118,112,125,117,101,77,132,128,45,86,48,60,148,185,225,159,219,214,219,214,103,175,180,175,182,179,177,217,222,221,219,212,118,122,124,158,160,106,133,129,50,64,79,47,80,134,133,129,112,107,93,101,149,208,206,206,98,144,142,130,119,131,127,124,129,170,165,65,32,187,152,172,158,156,178,157,157,172,128,122,127,130,126,127,133,133,121,122,114,137,137,78,78,69,71,79,84,97,165,137,115,197,189,171,166,159,167,163,183,179,99,67,84,97,104,101,70,73,105,72,68,86,92,96,114,121,111,127,120,124,126,123,117,102,84,109,133,140,23,55,65,56,139,191,225,163,219,215,217,223,158,178,178,169,173,175,165,218,222,220,217,212,118,127,116,171,166,88,131,115,80,84,53,51,71,110,110,163,138,92,124,144,176,208,206,200,87,142,125,116,99,120,120,118,124,151,163,56,22,143,166,184,181,168,169,119,120,148,124,101,118,121,124,64,132,99,106,93,69,117,117,78,78,65,79,73,80,160,163,121,196,197,148,144,129,113,108,102,124,123,98,108,97,110,119,108,80,87,91,104,113,112,110,119,130,155,131,113,131,141,135,176,213,214,217,192,136,135,25,27,50,56,138,193,211,171,210,219,224,218,170,170,176,168,171,182,171,218,220,217,216,213,127,140,116,170,166,70,127,127,115,112,56,41,43,59,47,152,143,88,125,126,196,205,204,204,84,129,129,102,94,154,104,99,108,144,157,48,25,182,185,184,182,186,181,184,181,174,180,166,141,144,140,160,160,160,128,105,65,110,110,77,77,75,72,80,82,134,134,95,128,142,132,168,105,107,86,80,93,126,139,133,138,139,140,124,106,84,101,132,135,124,204,196,208,215,209,163,210,213,211,216,218,219,222,181,129,128,19,41,42,32,92,174,211,193,209,219,220,217,187,164,170,171,167,181,175,215,218,216,218,215,135,147,125,152,163,68,132,114,107,84,46,34,33,39,34,147,145,114,114,130,183,207,205,201,114,101,143,88,85,105,91,99,108,137,139,60,32,193,192,185,179,178,181,180,181,182,186,185,185,185,184,182,177,178,180,181,174,149,149,98,98,83,94,85,75,151,168,98,115,122,123,201,153,118,135,122,125,135,157,157,154,153,157,139,133,117,163,134,150,136,136,150,117,207,169,116,192,218,221,221,215,222,217,114,134,135,43,37,36,26,114,185,196,209,199,220,220,222,212,151,175,169,168,178,183,209,214,220,217,225,132,143,133,159,165,66,124,47,53,40,39,30,36,30,33,108,103,100,86,91,157,204,203,199,90,67,83,78,73,83,92,100,99,128,132,61,136,190,180,174,175,181,181,177,182,186,181,183,182,180,186,183,180,178,177,182,185,181,181,131,131,78,136,82,79,101,130,87,90,101,119,203,205,128,159,154,156,145,160,162,161,160,153,186,151,144,79,154,151,133,142,111,138,111,106,130,115,163,223,203,138,219,221,91,104,104,67,45,41,34,94,174,150,194,187,210,209,205,205,150,170,171,165,172,181,172,212,215,216,209,132,144,139,162,126,61,72,30,37,53,26,28,29,112,106,122,89,101,68,95,195,201,204,205,196,89,103,103,106,95,60,111,106,113,104,101,190,181,187,180,173,178,175,182,183,180,183,175,177,181,176,179,181,181,177,173,172,171,171,130,130,129,155,85,82,84,98,111,111,102,109,202,205,133,174,167,173,165,159,148,151,159,156,165,191,135,197,154,160,150,165,117,92,91,89,167,108,102,98,123,98,204,220,93,179,155,154,86,89,48,185,193,169,207,187,210,213,205,198,155,183,197,198,199,185,155,204,206,204,203,141,135,78,106,125,118,33,30,107,48,45,79,64,125,164,149,80,51,28,102,108,208,206,201,204,107,93,77,122,71,35,78,106,111,118,175,181,179,182,182,161,171,177,175,173,176,179,176,184,176,179,178,178,179,179,177,176,178,178,162,162,140,132,99,103,87,100,118,112,122,109,204,207,165,167,175,165,165,147,147,146,154,163,157,209,117,162,138,127,134,158,152,144,141,87,106,122,122,110,95,95,202,202,104,167,156,160,172,132,153,193,189,181,197,163,215,215,219,209,186,195,197,199,199,199,161,215,214,212,211,182,134,136,129,141,122,94,78,119,30,150,131,191,157,178,129,103,102,84,94,111,131,203,205,200,82,47,89,154,98,57,86,114,136,142,165,178,173,183,182,114,153,161,172,166,170,176,174,176,181,173,173,178,180,175,173,175,175,175,111,111,106,109,115,118,96,152,117,114,126,117,192,200,176,155,173,163,161,147,150,149,165,165,168,157,132,160,169,208,215,223,213,217,195,211,109,101,123,107,97,93,111,123,108,162,152,155,155,137,149,192,193,167,195,176,217,214,220,216,217,186,192,191,195,192,173,208,216,219,209,171,124,127,130,128,159,144,149,157,148,154,129,136,150,156,133,62,128,71,100,151,152,205,201,199,88,51,69,76,68,53,47,119,106,174,137,162,162,180,170,111,139,156,167,161,165,172,169,167,174,174,172,178,182,180,181,182,176,176,119,119,110,101,104,106,104,137,119,111,99,117,190,197,186,159,160,163,147,152,159,165,167,174,173,169,147,146,141,166,161,155,152,151,140,176,164,152,124,137,182,208,97,126,119,150,155,146,143,124,146,188,195,163,184,185,217,219,217,219,217,148,180,183,190,190,188,196,215,215,214,144,116,137,125,131,128,89,110,160,154,142,135,123,147,153,168,167,146,30,136,163,139,207,197,200,168,37,174,111,150,166,187,79,130,193,172,139,145,181,183,122,165,173,165,149,158,164,162,164,157,164,165,170,175,178,182,182,178,178,139,139,127,122,105,110,105,121,116,118,107,114,176,203,199,163,161,159,166,175,163,164,173,197,170,149,137,178,196,152,161,145,216,119,209,140,116,216,213,169,124,201,106,124,106,148,129,118,108,131,135,186,189,147,179,189,214,213,201,215,215,151,174,184,193,197,187,189,215,212,215,145,120,121,128,111,108,82,141,139,154,149,104,138,153,151,174,139,130,41,148,159,201,190,192,193,116,34,178,186,181,178,135,38,35,177,196,185,202,181,178,151,147,172,167,121,143,157,157,147,138,147,159,164,167,174,171,169,180,180,150,150,134,157,114,120,107,107,112,112,114,109,153,201,200,168,165,162,175,162,161,167,198,213,200,177,206,218,208,203,165,200,214,189,216,208,206,224,222,216,187,144,114,119,107,146,139,157,127,126,129,183,175,135,151,202,215,217,180,189,209,189,177,179,183,191,201,175,215,216,212,125,131,137,118,106,102,69,75,111,153,153,128,127,113,127,145,145,177,161,134,104,164,73,191,133,65,131,189,182,185,187,150,143,71,68,193,200,196,198,173,130,143,166,150,84,137,148,162,138,103,144,150,139,143,169,171,166,183,183,130,130,142,122,155,103,122,136,125,103,114,112,189,196,198,177,169,161,177,177,196,198,195,196,199,201,201,200,195,200,198,210,206,209,208,215,211,211,214,211,221,219,136,97,106,152,151,150,108,112,112,158,172,124,147,211,207,160,161,141,186,172,105,176,176,189,202,170,207,218,217,144,127,123,90,104,73,46,73,129,132,122,124,110,86,96,80,103,119,131,118,76,62,62,61,137,151,157,183,176,185,171,178,174,55,65,62,64,77,124,196,196,187,175,199,99,150,141,158,150,99,132,152,140,177,177,190,178,145,145,149,149,116,115,143,115,123,145,118,122,108,117,181,196,201,198,190,199,199,201,195,197,190,190,200,199,195,200,206,207,209,207,208,209,211,200,211,214,212,210,217,219,218,208,98,124,137,135,101,101,87,174,184,136,190,204,190,156,146,123,128,107,73,163,177,183,193,181,194,214,215,152,119,109,98,66,39,89,81,124,123,120,102,98,81,106,106,128,110,124,87,83,61,98,107,154,172,177,184,184,183,180,156,176,113,59,62,65,63,62,63,174,196,193,196,122,133,128,146,146,73,106,155,151,140,170,148,163,144,144,145,145,150,145,108,106,114,138,130,151,130,171,195,197,198,196,194,194,193,194,202,203,184,188,191,193,187,192,199,198,206,209,198,205,198,195,196,203,210,208,207,213,223,215,90,90,95,111,72,89,118,184,185,140,186,185,146,143,110,54,57,69,58,61,110,176,180,183,180,219,211,160,116,74,81,93,100,120,94,92,100,100,83,80,89,103,123,136,130,126,126,129,91,115,137,128,158,158,166,170,170,163,190,190,118,61,66,70,61,63,64,69,141,199,197,193,99,111,134,138,124,137,130,165,126,155,161,164,178,178,154,154,156,154,119,115,147,192,197,207,203,205,201,212,206,210,197,192,202,177,177,176,114,123,130,96,92,187,168,179,126,118,175,172,185,209,205,213,202,211,213,203,118,125,119,74,117,130,95,91,101,83,156,102,164,189,114,99,64,54,34,110,41,40,32,172,189,175,169,219,208,169,92,59,73,115,128,111,78,76,93,76,85,84,74,79,98,95,120,93,126,93,88,95,101,197,128,158,153,120,174,166,157,153,86,45,47,53,62,71,65,56,65,69,68,106,178,156,87,161,93,136,119,192,198,183,189,182,193,193,184,184,187,192,200,201,203,206,205,203,206,210,207,206,207,198,147,137,167,197,182,207,135,87,99,111,131,108,103,114,97,116,99,108,94,121,110,131,162,193,195,104,107,97,104,69,127,127,94,104,211,197,193,142,144,133,67,47,47,174,99,103,103,88,73,178,163,185,176,193,208,160,137,160,183,193,173,183,133,100,77,85,82,122,105,86,113,167,171,189,188,168,162,167,173,181,172,177,166,167,166,165,168,147,56,35,45,37,39,41,58,53,73,70,74,73,57,64,177,196,189,189,200,195,190,201,196,162,190,190,191,191,195,194,202,203,202,204,205,207,205,209,209,207,192,162,161,198,212,214,213,208,117,216,212,154,199,184,94,101,102,96,165,138,134,146,149,141,150,118,16,64,76,39,83,62,51,114,95,114,148,138,191,127,135,58,48,22,79,108,104,147,123,166,176,178,204,205,194,140,127,52,203,207,177,200,193,53,127,124,113,123,115,120,133,126,170,183,178,181,178,177,180,175,179,181,175,174,167,171,168,176,164,162,148,137,113,130,115,100,111,54,64,61,85,135,112,179,177,180,154,169,201,201,186,197,197,135,188,188,194,194,194,194,199,202,201,203,208,202,212,206,205,208,210,210,209,209,208,215,214,211,211,217,214,215,214,214,214,191,91,103,138,147,157,146,145,139,144,128,126,108,109,89,93,109,41,100,91,131,147,125,215,105,165,50,148,184,179,141,182,129,137,48,167,166,147,154,153,145,126,60,165,79,66,91,198,57,75,128,128,123,85,50,88,194,54,91,177,185,180,189,187,185,186,179,180,175,182,173,177,173,176,182,168,172,169,158,152,89,78,80,68,103,106,152,121,140,165,118,127,143,165,161,162,168,162,130,177,177,196,196,191,197,200,200,203,204,205,207,204,205,207,207,206,208,209,209,210,209,211,211,212,211,215,211,212,211,210,213,201,197,198,191,165,164,146,89,131,146,105,117,136,122,161,155,161,156,151,125,119,131,82,84,103,32,146,132,87,89,87,112,172,72,171,108,58,99,172,168,170,171,132,164,168,187,193,178,177,99,152,123,176,175,149,180,155,163,180,185,190,187,185,185,183,181,185,180,176,180,179,181,176,180,171,143,168,161,153,119,114,91,74,103,111,124,134,150,174,120,135,166,147,118,144,170,138,123,100,100,195,195,196,197,199,201,202,204,205,204,203,207,205,205,207,206,209,210,207,214,207,209,210,212,200,176,205,206,204,194,211,197,217,218,203,196,183,142,138,175,207,210,76,86,169,196,182,180,186,183,171,138,153,160,161,158,143,115,91,104,77,95,127,95,71,186,160,171,183,182,181,179,172,176,177,180,172,162,169,164,166,162,164,168,169,162,175,172,179,181,180,175,175,177,177,175,172,177,177,178,179,173,175,180,177,175,146,116,161,114,110,64,76,110,113,118,128,133,139,132,135,115,105,130,126,154,84,92,104,104,196,196,195,195,198,201,203,204,205,203,201,205,205,203,203,205,213,211,208,211,212,213,201,154,142,150,159,180,194,189,157,151,161,201,180,149,163,112,189,208,209,211,106,114,115,205,200,196,166,137,129,131,154,167,160,159,155,158,167,162,167,141,119,150,130,160,168,178,167,174,181,176,180,183,180,182,180,176,179,176,177,179,181,182,175,179,178,179,177,169,159,149,160,160,168,165,179,175,180,181,176,175,176,169,176,174,135,127,152,108,104,98,107,115,116,117,98,135,69,115,130,101,97,118,113,131,70,99,105,105,193,193,194,197,201,201,199,199,200,205,202,203,204,205,205,203,205,210,206,202,187,156,164,163,152,158,147,126,173,168,129,73,117,208,208,206,211,216,132,212,189,212,210,198,205,201,204,203,173,102,118,124,149,163,170,163,168,164,168,165,171,176,172,177,175,177,183,183,182,181,174,182,184,178,180,185,183,182,182,184,182,157,175,167,170,166,165,163,160,157,160,173,171,176,176,169,170,174,176,176,175,182,183,177,178,172,147,129,119,125,101,81,76,115,108,75,52,69,52,59,108,104,116,115,111,106,81,82,98,98,196,196,196,197,199,200,200,200,202,198,202,204,200,197,200,203,204,202,190,167,161,170,167,162,160,145,150,103,164,73,110,144,120,204,209,213,217,212,77,195,182,187,195,203,208,211,199,198,82,89,123,150,141,159,161,162,163,163,165,163,167,164,164,173,178,190,185,194,190,182,182,182,173,176,181,184,180,182,183,186,177,146,152,148,152,156,148,151,165,164,172,175,179,174,177,173,178,178,179,168,171,171,173,171,174,109,149,122,98,101,37,28,47,92,77,38,60,68,44,56,102,106,64,96,96,92,99,88,99,99,197,197,196,196,198,200,200,199,198,202,198,196,199,197,193,194,197,186,163,170,174,178,165,152,150,139,141,117,134,140,156,52,38,70,197,209,216,190,73,181,180,175,161,156,170,177,193,194,197,138,84,192,81,84,138,156,155,157,161,170,164,160,166,165,174,167,179,179,185,189,182,187,175,171,174,177,176,179,175,165,145,143,142,138,135,145,165,159,172,171,174,175,177,174,179,170,172,176,176,167,166,171,172,162,126,75,109,44,65,122,51,34,32,51,39,32,49,66,43,48,60,53,66,95,84,86,83,85,93,93,192,192,196,199,199,199,200,201,202,190,197,197,195,198,200,188,166,176,172,172,168,161,158,155,151,144,79,115,33,92,142,42,28,81,189,129,164,60,12,141,166,156,153,151,151,154,171,180,161,164,157,179,178,144,122,141,115,124,131,154,171,169,163,167,168,170,166,167,169,173,164,159,163,166,165,169,171,171,165,155,145,126,166,154,167,150,161,171,165,163,168,170,169,174,171,173,169,173,180,172,159,109,146,125,70,65,54,60,65,62,52,19,48,30,121,43,44,45,42,43,99,48,54,72,81,73,87,67,77,77,193,193,197,198,197,197,200,201,198,201,191,180,180,175,165,167,172,175,180,170,171,164,155,152,146,148,130,137,148,165,168,137,131,150,175,158,138,121,145,162,172,162,154,170,162,157,167,167,169,165,170,156,148,159,187,200,164,148,126,112,128,162,165,165,170,170,165,163,163,161,158,166,157,154,152,155,153,148,152,156,165,170,163,162,153,144,156,160,168,163,149,170,168,159,169,137,161,126,176,74,100,76,83,46,59,64,65,58,59,67,29,36,26,28,28,33,38,45,28,33,37,46,33,47,71,69,78,57,56,56,193,193,195,197,199,201,196,177,157,149,153,155,164,169,171,178,180,182,178,177,168,157,152,150,149,130,27,58,149,169,166,158,135,147,166,153,159,162,151,169,149,143,163,169,170,173,175,183,185,181,166,168,156,156,164,172,179,181,177,176,154,153,169,183,171,164,161,169,164,157,158,162,154,149,153,160,156,146,151,149,157,168,166,164,158,143,163,167,167,151,157,156,162,166,167,169,166,173,174,166,171,122,153,153,83,54,64,45,51,48,59,63,104,48,21,14,28,20,15,35,29,60,33,30,52,58,49,49,103,103,196,196,191,174,184,167,132,134,151,156,153,163,168,175,179,186,185,180,180,176,173,164,150,145,156,136,146,149,156,168,175,162,148,135,146,145,160,162,159,161,162,165,162,175,169,167,175,181,179,183,175,166,161,162,156,166,163,167,179,181,181,109,136,167,186,184,164,159,163,145,136,144,158,149,157,155,157,156,158,158,170,173,173,177,178,170,166,167,165,165,165,161,167,173,165,168,182,166,162,181,171,181,175,170,170,168,171,168,135,73,75,62,47,60,24,19,25,24,32,37,14,24,33,26,36,37,60,46,80,80,164,164,157,146,125,130,129,145,153,156,156,166,169,178,180,180,183,183,180,180,166,159,155,152,156,159,160,148,147,167,171,169,160,129,147,151,162,162,162,168,167,167,174,170,175,163,164,180,175,178,180,165,167,161,167,160,159,153,161,184,189,182,176,143,132,123,189,186,166,131,102,124,123,150,149,154,160,168,162,170,172,175,179,182,181,178,172,169,168,163,164,172,170,166,169,163,165,161,155,171,173,175,178,171,169,166,165,164,154,168,158,162,125,158,163,156,153,145,135,157,142,142,130,126,120,86,28,29,26,26,153,153,138,128,122,143,155,155,154,155,162,167,171,179,177,179,185,182,178,173,169,166,161,161,153,152,165,165,157,170,176,167,159,145,149,150,167,170,162,165,169,172,172,173,170,173,154,163,180,170,177,169,163,171,166,160,166,164,145,142,186,190,189,186,90,95,94,93,73,91,96,82,119,134,146,160,158,162,163,165,176,176,183,183,181,181,175,166,166,160,167,166,164,163,168,165,167,164,162,165,175,175,174,171,163,165,152,148,135,134,150,159,161,160,147,156,151,142,159,156,150,140,150,159,144,151,147,138,103,103,135,135,139,138,142,146,151,155,160,158,169,168,177,183,179,184,180,172,165,168,170,165,152,152,145,150,153,173,139,165,172,172,159,139,159,162,164,164,159,160,160,153,165,173,183,174,166,157,161,178,177,168,168,163,165,171,168,168,166,149,154,188,190,195,186,158,116,92,104,92,140,192,177,139,131,135,155,150,160,164,173,174,178,178,178,179,176,169,167,170,165,167,170,163,164,170,169,167,168,156,187,186,176,161,146,136,134,126,119,120,126,133,152,190,130,143,137,151,160,157,150,151,155,146,146,132,135,121,75,75,153,153,148,146,147,152,151,154,158,156,167,172,172,162,158,163,158,152,147,149,160,152,155,147,148,152,160,180,165,162,167,157,152,135,160,162,154,152,142,134,132,135,144,160,174,177,178,143,167,172,175,160,168,172,172,171,168,169,175,165,162,157,184,187,192,195,198,187,121,161,163,131,144,144,150,183,123,140,156,157,154,154,150,151,158,165,170,168,161,165,162,165,163,164,164,168,174,175,175,160,186,188,173,144,132,136,117,129,126,124,128,132,135,126,113,150,118,110,125,140,151,144,142,131,131,116,125,128,122,122,164,164,154,155,156,152,157,148,155,161,160,164,157,146,151,149,147,141,144,135,142,145,141,148,146,147,158,171,175,160,137,134,135,157,158,154,153,148,123,113,119,132,145,147,153,155,160,154,145,158,179,168,155,171,181,182,170,165,174,183,174,172,164,153,167,185,192,195,198,185,152,148,128,103,106,171,111,128,136,146,147,141,142,147,146,137,135,141,142,147,159,159,164,166,161,164,161,167,171,108,163,112,194,127,133,131,121,120,124,128,129,125,123,129,118,123,119,102,117,129,124,127,126,139,181,184,188,191,193,193,165,165,165,162,161,151,162,150,149,157,148,139,142,148,157,151,143,144,132,95,123,127,134,132,146,146,158,151,177,173,159,144,140,152,149,150,141,126,109,110,110,105,119,116,128,130,139,126,123,165,166,164,154,158,169,177,178,156,180,178,178,180,176,158,167,170,190,197,200,199,175,165,160,115,113,99,89,99,116,131,144,148,142,141,145,149,150,149,148,149,145,144,153,146,151,156,167,166,169,135,78,109,111,94,108,97,92,119,112,114,123,136,146,150,128,138,122,108,113,123,122,125,122,126,134,138,144,126,138,138,175,175,169,166,170,163,142,138,133,148,158,144,156,156,146,149,143,128,45,23,40,120,126,119,136,138,148,137,145,166,162,152,145,151,147,150,136,119,115,115,95,107,117,119,117,120,121,120,100,128,158,169,118,160,165,161,155,169,176,175,181,177,173,166,168,181,185,167,156,163,165,177,184,181,169,151,117,110,114,119,127,127,127,128,134,142,143,143,149,151,145,148,143,149,141,82,145,159,146,125,92,125,110,105,104,114,130,139,148,159,152,165,157,155,141,136,142,140,118,111,115,122,119,126,135,138,133,146,134,134,179,179,172,168,163,138,144,143,155,166,164,145,158,155,144,143,137,28,16,25,73,123,122,122,142,150,152,146,145,154,162,152,148,150,148,147,132,115,118,116,110,111,114,120,120,119,118,131,111,93,129,159,136,158,167,170,173,170,183,182,178,176,167,147,180,185,184,173,162,161,162,161,198,205,171,142,116,125,122,134,118,120,111,118,123,140,122,125,132,140,142,136,148,146,141,123,72,71,85,119,124,123,130,131,138,136,150,145,154,158,163,166,162,158,159,151,157,149,135,124,115,105,114,116,120,122,132,144,138,138,163,163,149,132,123,139,136,152,164,169,156,127,139,144,144,141,127,48,99,129,126,115,120,126,141,148,139,152,150,146,160,149,153,154,155,141,116,124,131,130,130,121,125,111,110,108,118,126,121,121,105,128,150,160,159,160,162,172,180,172,180,179,163,118,184,177,183,167,160,157,157,161,157,160,176,168,140,121,133,139,129,107,103,111,116,128,120,113,119,123,120,126,125,107,95,99,97,85,82,79,83,71,77,74,111,148,159,157,156,158,167,159,160,154,142,142,151,138,124,114,126,110,117,114,108,100,113,107,135,135,161,161,132,125,136,145,142,138,160,150,131,129,118,123,132,135,125,116,117,124,118,124,134,152,147,140,142,157,162,143,83,60,104,140,147,105,128,149,148,139,107,119,127,110,103,106,109,59,89,120,134,162,158,161,163,170,164,170,167,178,173,167,160,150,160,162,160,144,138,133,135,160,160,159,157,150,162,175,176,145,127,109,113,105,108,111,109,101,111,111,113,121,100,88,87,88,99,101,112,109,89,79,85,81,96,82,151,156,157,159,159,155,161,158,150,121,116,100,108,115,100,99,96,101,100,105,108,97,107,107,144,144,129,142,139,147,152,143,141,128,130,129,92,113,114,130,130,114,122,128,146,125,140,149,160,144,142,163,165,160,158,60,119,164,89,82,82,128,150,149,78,126,132,136,141,139,124,55,52,106,148,162,164,164,167,164,166,162,170,161,140,142,151,160,169,156,104,116,142,146,138,128,123,88,99,129,152,151,159,144,124,116,129,124,110,99,103,109,106,113,108,115,115,106,103,104,103,109,116,115,122,108,103,94,88,89,92,151,161,155,135,122,133,149,155,150,118,96,80,94,99,94,90,96,87,99,95,96,96,96,144,144,148,145,143,136,131,119,113,106,101,104,86,120,116,104,159,140,122,150,131,86,80,86,79,68,72,168,171,121,153,137,162,164,155,66,86,82,129,157,99,120,185,167,186,155,150,70,41,152,160,166,155,166,159,164,170,169,167,135,123,133,127,170,164,164,117,98,124,127,131,127,66,84,93,117,74,68,71,112,119,105,140,137,129,120,109,102,108,120,132,111,113,114,110,108,101,104,110,109,113,119,108,109,73,71,83,114,122,115,91,98,114,119,122,135,139,101,77,88,96,97,85,101,106,92,100,98,90,90,142,142,138,132,125,124,127,120,108,101,89,95,108,103,138,129,141,135,128,147,71,72,71,72,78,78,67,167,170,130,89,101,160,162,164,153,157,87,74,149,158,92,155,167,174,88,51,150,163,153,163,154,159,153,140,143,152,151,142,116,121,128,125,160,161,143,142,102,90,110,128,116,109,108,105,100,100,116,137,123,93,84,84,124,134,134,128,123,113,110,103,110,119,115,109,112,190,190,159,105,110,111,113,112,78,77,68,112,110,98,92,75,80,94,99,90,83,116,75,76,63,94,73,76,98,91,99,103,91,91,133,133,128,123,144,133,134,102,96,110,123,145,153,134,150,104,121,121,146,163,151,144,139,109,133,149,83,167,174,165,83,86,88,107,160,173,169,168,92,83,149,93,108,176,185,133,14,172,163,160,139,138,131,131,117,97,125,116,73,78,73,99,106,104,113,120,132,111,98,84,114,121,123,114,95,100,109,102,109,137,147,191,128,58,101,123,130,140,132,120,116,108,114,110,112,111,124,178,173,171,177,172,146,129,68,79,84,120,119,117,88,90,60,73,73,73,74,105,79,69,69,86,72,71,117,168,172,171,156,156,101,101,141,141,135,130,120,122,129,152,147,153,157,168,161,103,113,153,154,140,133,146,127,109,103,129,105,140,131,115,80,84,85,82,81,127,165,143,61,35,94,88,89,116,134,135,133,140,123,124,134,92,94,90,87,92,73,100,102,99,96,85,86,78,85,79,82,94,112,78,100,107,114,104,101,100,101,154,160,167,151,113,125,130,86,86,77,114,145,144,142,133,117,114,108,108,168,172,163,173,167,166,171,172,92,90,112,110,105,106,105,107,116,74,76,70,97,93,71,70,72,95,89,136,171,172,162,168,159,159,118,118,140,139,132,135,133,131,153,154,134,136,145,175,157,91,112,101,84,91,86,81,88,94,107,82,104,119,123,114,81,82,80,90,53,70,158,135,85,81,94,70,88,101,87,86,117,105,109,109,85,100,92,68,75,93,83,92,116,75,55,111,78,70,56,100,80,78,71,78,69,98,107,105,98,103,91,134,145,162,160,161,146,101,102,110,84,75,65,109,155,149,136,123,122,111,131,150,171,172,169,178,172,147,118,102,121,141,123,113,108,104,96,99,83,93,112,103,99,68,93,90,145,178,172,175,169,162,157,157,132,132,141,137,134,131,134,136,133,130,120,109,111,144,120,103,98,100,94,95,97,102,95,106,102,86,102,99,98,92,84,83,78,90,93,99,100,87,63,95,86,88,82,100,95,62,85,122,109,108,81,85,94,98,75,87,89,91,95,89,97,110,107,104,98,91,89,83,66,70,63,40,67,105,99,94,104,107,156,163,157,169,154,148,127,98,108,88,59,90,81,122,148,142,136,127,130,136,135,145,146,159,169,111,111,118,109,169,171,153,144,114,99,97,79,104,98,100,100,88,96,84,94,133,156,168,159,157,158,158,133,133,146,139,137,130,124,134,144,154,156,124,124,128,133,129,136,134,123,124,105,101,103,75,92,87,89,90,103,95,80,72,81,92,92,99,100,99,61,89,75,92,80,97,99,89,74,108,119,99,86,83,84,92,71,81,88,93,92,71,81,93,108,103,71,75,77,77,86,101,88,54,22,67,103,106,90,71,100,92,103,104,97,93,93,93,90,65,73,72,53,35,54,105,136,135,129,126,134,132,137,137,150,77,91,108,103,179,179,181,178,141,134,155,115,108,90,89,96,113,96,85,79,90,81,84,143,159,154,154,165,165,167,160,166,166,160,153,147,142,135,140,133,131,133,139,134,140,139,138,93,108,106,72,84,89,84,83,89,93,86,81,87,96,91,92,89,100,93,69,81,78,84,84,97,104,80,99,111,100,78,88,94,87,80,72,94,92,83,63,11,48,91,94,20,36,69,46,104,102,15,102,63,101,91,94,108,45,88,89,93,100,99,101,99,94,96,99,88,73,65,38,25,38,48,76,77,87,96,100,94,117,116,74,77,84,79,128,152,174,180,147,141,168,171,172,126,90,81,108,120,123,106,98,111,97,88,79,117,117,172,172,181,168,154,149,139,117,111,112,131,128,139,131,140,128,115,89,83,85,85,102,100,61,76,74,81,89,92,97,97,89,87,81,82,84,101,96,93,57,63,68,64,68,77,72,76,68,92,96,71,61,87,83,65,68,85,56,69,70,73,78,90,95,87,97,106,93,113,113,108,121,123,111,115,121,98,78,90,88,90,99,96,97,88,87,89,82,82,88,61,53,26,45,25,27,36,54,74,81,66,111,107,67,90,79,74,67,96,112,110,110,171,177,183,184,187,180,153,159,125,114,120,113,120,124,116,109,94,94,151,151,140,133,124,109,112,109,102,105,99,95,113,98,96,93,93,97,95,87,80,91,83,83,71,71,77,79,84,79,76,72,82,65,81,90,90,100,102,63,64,65,59,66,73,78,75,70,79,101,73,69,67,75,58,61,92,50,84,77,81,91,94,106,96,104,111,122,119,125,109,117,115,115,108,110,78,73,74,84,90,89,91,91,89,82,82,69,80,90,94,101,54,51,55,52,44,39,39,27,36,78,107,71,80,88,93,90,88,84,79,76,85,135,149,166,178,175,182,198,196,191,175,153,123,109,124,125,109,109,125,125,120,112,114,110,104,99,103,96,102,100,87,85,93,87,91,88,85,89,83,80,81,72,73,77,78,72,70,68,67,64,65,67,76,80,90,105,102,93,82,77,67,90,80,88,87,81,60,62,54,69,81,101,61,63,86,84,79,76,82,89,99,103,100,60,63,123,131,124,116,111,114,109,104,96,60,55,53,61,67,65,68,69,77,65,56,56,76,94,103,110,109,93,83,75,76,78,66,74,59,37,36,55,61,75,84,96,97,109,99,98,89,98,134,133,127,137,165,173,183,194,197,200,196,189,178,122,112,112,128,128,131,118,124,127,112,96,90,89,89,85,80,82,83,80,86,82,88,86,79,86,80,77,81,73,73,71,64,67,57,62,63,62,67,73,81,91,94,89,93,93,98,103,108,126,127,127,117,107,96,85,87,104,64,78,85,87,83,73,77,106,97,106,110,98,99,100,125,119,120,115,108,102,86,95,99,100,87,85,82,80,66,67,64,60,63,62,61,66,73,80,97,99,102,103,104,88,84,88,81,87,61,60,89,67,83,95,109,110,119,135,130,125,116,136,135,155,181,183,181,179,181,185,194,192,193,189,187,187,128,128,131,118,124,127,112,96,90,89,89,85,80,82,83,80,86,82,88,86,79,86,80,77,81,73,73,71,64,67,57,62,63,62,67,73,81,91,94,89,93,93,98,103,108,126,127,127,117,107,96,85,87,104,64,78,85,87,83,73,77,106,97,106,110,98,99,100,125,119,120,115,108,102,86,95,99,100,87,85,82,80,66,67,64,60,63,62,61,66,73,80,97,99,102,103,104,88,84,88,81,87,61,60,89,67,83,95,109,110,119,135,130,125,116,136,135,155,181,183,181,179,181,185,194,192,193,189,187,187};
    


module controller_tb();
    logic clk;
    logic reset;
    logic done;
    logic stall;
    logic [12:0] address_read;
    logic [12:0] address_write;
    logic [7:0]data_in;
    logic [7:0]temp_out[8:0];
    logic signed [7:0] fil [0:2][0:2]='{'{0,-1,0}, {-1,5,-1}, {0,-1,0}};
   


    always@(negedge clk)begin
    
        data_in=arar[address_read];
    
    end

    Top_module mod(fil,stall,Recieve, RxD, TxD, clk, reset, Transmitt, done, done_out,data_in,address_read);
     
     initial begin
     clk=0;
     forever begin
     clk=~clk; #5;
     end
     end
     
     initial begin
     reset=1;
     stall=1;
     #15;
     stall=0;
     reset=0;
     done=1;
     #50;
     end
     
 endmodule